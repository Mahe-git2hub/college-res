module _42encoder_tb;
reg a3,a2,a1,a0;
wire f1,f0;
fourtwoencoder my_gate(a3,a2,a1,a0,f1,f0);
initial 
begin 
$monitor("a3=%b a2=%b a1=%b a0=%b f1=%b f0=%b",a3,a2,a1,a0,f1,f0);
a3=1'b0;
a2=1'b0;
a1=1'b0;
a0=1'b0;
#10;
a3=1'b0;
a2=1'b0;
a1=1'b0;
a0=1'b1;
#10;
a3=1'b0;
a2=1'b0;
a1=1'b1;
a0=1'b0;
#10;
a3=1'b0;
a2=1'b0;
a1=1'b1;
a0=1'b1;
#10;
a3=1'b0;
a2=1'b1;
a1=1'b0;
a0=1'b0;
#10;
a3=1'b0;
a2=1'b1;
a1=1'b0;
a0=1'b1;
#10;
a3=1'b0;
a2=1'b1;
a1=1'b1;
a0=1'b0;
#10;
a3=1'b0;
a2=1'b1;
a1=1'b1;
a0=1'b1;
#10;
a3=1'b1;
a2=1'b0;
a1=1'b0;
a0=1'b0;
#10;
a3=1'b1;
a2=1'b0;
a1=1'b0;
a0=1'b1;
#10;
a3=1'b1;
a2=1'b0;
a1=1'b1;
a0=1'b0;
#10;
a3=1'b1;
a2=1'b0;
a1=1'b1;
a0=1'b1;
#10;
a3=1'b1;
a2=1'b1;
a1=1'b0;
a0=1'b0;
#10;
a3=1'b1;
a2=1'b1;
a1=1'b0;
a0=1'b1;
#10;
a3=1'b1;
a2=1'b1;
a1=1'b1;
a0=1'b0;
#10;
a3=1'b1;
a2=1'b1;
a1=1'b1;
a0=1'b1;
end
endmodule